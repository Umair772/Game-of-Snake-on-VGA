//Umair Liaqat
//12/6/2019
//Umair and Abdiasis
module generateAppleCoordinates (CLOCK_50,x,y,start,reset,good_collision,apple);
	//Declaring input and output logics
	input logic CLOCK_50,reset,good_collision,start;
	output logic [7:0]apple; //Outputs a 8-bit apple location
	logic [7:0]appleX; //X-coordinate for the apple
   logic [7:0]appleY; //Y-coordinate for the apple
   logic [9:0]appX;   //random values generated by the LFSR
   logic [9:0]appY;   //random values generated by the LFSR
	logic [7:0]inX,inY; //Makes the pixel on the screen
	input logic [9:0]x; //X pixel
	input logic [8:0]y; //Y pixel
   
	//10-bit LFSRs which outputs a random value
	LFSR #(.n(10)) randX (.clk(CLOCK_50),.reset(reset),.start(start),.out(appX));
	LFSR #(.n(10)) randY (.clk(CLOCK_50),.reset(reset),.start(start),.out(appY));
	
   //flip flop which is reponsible for reset and starting the game. To make sure the apple is generated within the borders.
	always_ff @(posedge CLOCK_50) begin
		if (reset || ~start) begin
			appleX <= 300;
			appleY <= 350;
		end
		else begin
		   if (good_collision) begin
			   if((appX<10) || (appX>630) || (appY<10) || (appY>470)) begin
				   appleX <= 40;
				   appleY <= 30;
			   end
			   else begin
					appleX <= appX;
					appleY <= appY;
		    end
		 end
	  end
	end
	
  //Using a flip flop to make a pixel on the screen by using the coordinates provided by the VGA driver.	
  always @(posedge CLOCK_50)
	  begin
		 inX <= (x > (appleX - 10) && x < (appleX + 10));
		 inY <= (y > (appleY - 10) && y < (appleY + 10));
	  end
	  
	assign apple = inX && inY;
	  

endmodule

//Simulating in modelsim
module generateAppleCoordinates_testbench();

   logic CLOCK_50,reset,good_collision,gameOver;
	logic [9:0]x,y;
   logic [9:0]appleX;
   logic [9:0]appleY;
	logic [9:0]appX;
	logic [9:0]appY;
	logic apple,r,g,b;
	logic inX,inY;
   logic [7:0] VGA_R,VGA_G,VGA_B;
   logic VGA_BLANK_N;
   logic VGA_CLK;
   logic VGA_HS;
   logic VGA_SYNC_N;
   logic VGA_VS;
	
	
	generateAppleCoordinates dut (.CLOCK_50,.reset,.good_collision,.gameOver,.apple,.VGA_R,.VGA_G,.VGA_B,.VGA_CLK,.VGA_BLANK_N,.VGA_HS,.VGA_SYNC_N,.VGA_VS);
	
	
	parameter CLOCK_PERIOD = 100;
	initial CLOCK_50 = 1;
	always begin
	    #(CLOCK_PERIOD/2);
		 CLOCK_50 = ~CLOCK_50;
	end
	
	initial begin
	reset <= 1;       @(posedge CLOCK_50);
	reset <= 0;					@(posedge CLOCK_50);
	good_collision <= 1; gameOver <= 0; 						@(posedge CLOCK_50);
	good_collision <= 0; 						@(posedge CLOCK_50);
							@(posedge CLOCK_50);
							@(posedge CLOCK_50);
							@(posedge CLOCK_50);
							@(posedge CLOCK_50);
							@(posedge CLOCK_50);
							@(posedge CLOCK_50);
							@(posedge CLOCK_50);
							@(posedge CLOCK_50);
  good_collision <= 1;							@(posedge CLOCK_50);
  good_collision <= 0; 							@(posedge CLOCK_50);
							@(posedge CLOCK_50);
							@(posedge CLOCK_50);
							@(posedge CLOCK_50);
							@(posedge CLOCK_50);
							@(posedge CLOCK_50);
							@(posedge CLOCK_50);
							@(posedge CLOCK_50);
							@(posedge CLOCK_50);
							@(posedge CLOCK_50);
							@(posedge CLOCK_50);
							@(posedge CLOCK_50);
  $stop();
  end
 endmodule

			
	
	